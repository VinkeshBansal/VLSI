magic
tech scmos
timestamp 1669566576
<< error_s >>
rect -953 769 -952 774
rect -1175 684 -1174 689
rect -952 394 -951 399
rect -1174 309 -1173 314
rect -911 306 -905 307
rect -952 16 -951 21
rect -1174 -69 -1173 -64
rect 140 -90 141 -85
rect -82 -175 -81 -170
rect -1345 -420 -1344 -415
rect 141 -465 142 -460
rect -81 -550 -80 -545
rect 182 -553 188 -552
rect 141 -843 142 -838
rect -81 -928 -80 -923
rect 1246 -949 1247 -944
rect -252 -1279 -251 -1274
rect 1247 -1324 1248 -1319
rect 1288 -1412 1294 -1411
rect 1247 -1702 1248 -1697
rect 854 -2138 855 -2133
<< metal1 >>
rect -1719 873 -1551 882
rect -1719 600 -1551 604
rect -838 590 -772 594
rect -621 591 -617 623
rect -838 504 -832 590
rect -706 587 -617 591
rect -706 580 -646 584
rect -841 496 -832 504
rect -821 504 -772 508
rect -621 505 -617 587
rect -821 466 -815 504
rect -706 501 -617 505
rect -706 494 -646 498
rect -841 458 -815 466
rect -841 429 -826 437
rect -831 422 -826 429
rect -831 418 -772 422
rect -621 419 -617 501
rect -706 415 -617 419
rect -706 408 -646 412
rect -841 395 -828 403
rect -835 336 -828 395
rect -835 332 -772 336
rect -621 333 -617 415
rect -706 329 -617 333
rect -706 322 -646 326
rect -1719 225 -1551 229
rect -840 24 -458 34
rect -462 14 -458 24
rect -841 1 -470 12
rect -840 -41 -519 -31
rect -840 -64 -580 -54
rect -1719 -153 -1551 -149
rect -1719 -504 -1551 -500
rect -590 -1008 -580 -64
rect -528 -630 -519 -41
rect -481 -255 -471 1
rect -481 -259 -458 -255
rect 255 -269 321 -265
rect 472 -268 476 -236
rect 255 -355 261 -269
rect 387 -272 476 -268
rect 387 -279 447 -275
rect 252 -363 261 -355
rect 272 -355 321 -351
rect 472 -354 476 -272
rect 272 -393 278 -355
rect 387 -358 476 -354
rect 387 -365 447 -361
rect 252 -401 278 -393
rect 252 -430 267 -422
rect 262 -437 267 -430
rect 262 -441 321 -437
rect 472 -440 476 -358
rect 387 -444 476 -440
rect 387 -451 447 -447
rect 252 -464 265 -456
rect 258 -523 265 -464
rect 258 -527 321 -523
rect 472 -526 476 -444
rect 387 -530 476 -526
rect 387 -537 447 -533
rect -528 -634 -458 -630
rect 253 -835 647 -825
rect 640 -837 647 -835
rect 640 -844 648 -837
rect 252 -858 623 -847
rect 253 -900 574 -890
rect 253 -923 513 -913
rect -590 -1012 -458 -1008
rect -1719 -1359 -1706 -1358
rect -1719 -1363 -458 -1359
rect 503 -1867 513 -923
rect 565 -1489 574 -900
rect 612 -1114 622 -858
rect 612 -1118 648 -1114
rect 1361 -1128 1427 -1124
rect 1578 -1127 1582 -1095
rect 1361 -1214 1367 -1128
rect 1493 -1131 1582 -1127
rect 1493 -1138 1553 -1134
rect 1358 -1222 1367 -1214
rect 1378 -1214 1427 -1210
rect 1578 -1213 1582 -1131
rect 1378 -1252 1384 -1214
rect 1493 -1217 1582 -1213
rect 1493 -1224 1553 -1220
rect 1358 -1260 1384 -1252
rect 1358 -1289 1373 -1281
rect 1368 -1296 1373 -1289
rect 1368 -1300 1427 -1296
rect 1578 -1299 1582 -1217
rect 1493 -1303 1582 -1299
rect 1493 -1310 1553 -1306
rect 1358 -1323 1371 -1315
rect 1364 -1382 1371 -1323
rect 1364 -1386 1427 -1382
rect 1578 -1385 1582 -1303
rect 1493 -1389 1582 -1385
rect 1493 -1396 1553 -1392
rect 565 -1493 648 -1489
rect 1359 -1694 1366 -1641
rect 1377 -1687 1432 -1683
rect 1582 -1686 1586 -1637
rect 1377 -1707 1382 -1687
rect 1498 -1690 1586 -1686
rect 1498 -1697 1558 -1693
rect 1359 -1717 1382 -1707
rect 1359 -1759 1386 -1749
rect 1381 -1769 1386 -1759
rect 1359 -1855 1365 -1772
rect 1381 -1773 1432 -1769
rect 1582 -1772 1586 -1690
rect 1498 -1776 1586 -1772
rect 1497 -1783 1557 -1779
rect 1359 -1859 1432 -1855
rect 1582 -1858 1586 -1776
rect 1498 -1862 1586 -1858
rect 503 -1871 648 -1867
rect 1498 -1869 1558 -1865
rect -1719 -2218 -677 -2217
rect -1719 -2221 648 -2218
rect -717 -2222 648 -2221
rect -1719 -2315 1432 -2311
rect 1582 -2314 1586 -1862
rect 1498 -2318 1586 -2314
rect 1498 -2325 1558 -2321
use Adder_4  Adder_4_2
timestamp 1669566576
transform 0 1 -1458 -1 0 499
box -382 -93 1069 618
use AND  AND_11
timestamp 1669566576
transform -1 0 -706 0 -1 621
box 0 0 66 83
use AND  AND_12
timestamp 1669566576
transform -1 0 -706 0 -1 535
box 0 0 66 83
use AND  AND_13
timestamp 1669566576
transform -1 0 -706 0 -1 449
box 0 0 66 83
use AND  AND_14
timestamp 1669566576
transform -1 0 -706 0 -1 363
box 0 0 66 83
use Adder_4  Adder_4_1
timestamp 1669566576
transform 0 1 -365 -1 0 -360
box -382 -93 1069 618
use AND  AND_9
timestamp 1669566576
transform -1 0 387 0 -1 -238
box 0 0 66 83
use AND  AND_10
timestamp 1669566576
transform -1 0 387 0 -1 -324
box 0 0 66 83
use AND  AND_8
timestamp 1669566576
transform -1 0 387 0 -1 -410
box 0 0 66 83
use AND  AND_3
timestamp 1669566576
transform -1 0 387 0 -1 -496
box 0 0 66 83
use Adder_4  Adder_4_0
timestamp 1669566576
transform 0 1 741 -1 0 -1219
box -382 -93 1069 618
use AND  AND_5
timestamp 1669566576
transform -1 0 1493 0 -1 -1097
box 0 0 66 83
use AND  AND_4
timestamp 1669566576
transform -1 0 1493 0 -1 -1183
box 0 0 66 83
use AND  AND_6
timestamp 1669566576
transform -1 0 1493 0 -1 -1269
box 0 0 66 83
use AND  AND_7
timestamp 1669566576
transform -1 0 1493 0 -1 -1355
box 0 0 66 83
use AND  AND_2
timestamp 1669566576
transform -1 0 1498 0 -1 -1656
box 0 0 66 83
use AND  AND_1
timestamp 1669566576
transform -1 0 1498 0 -1 -1742
box 0 0 66 83
use AND  AND_0
timestamp 1669566576
transform -1 0 1498 0 -1 -1828
box 0 0 66 83
use AND  AND_15
timestamp 1669566576
transform -1 0 1498 0 -1 -2284
box 0 0 66 83
<< labels >>
rlabel metal1 -1713 -2315 -1713 -2311 3 P0
rlabel metal1 -1714 -2221 -1714 -2217 3 P1
rlabel metal1 -1713 -1362 -1713 -1358 3 P2
rlabel metal1 -1714 -504 -1714 -500 3 P3
rlabel metal1 -1714 -153 -1714 -149 3 P4
rlabel metal1 -1712 225 -1712 229 3 P5
rlabel metal1 -1714 600 -1714 604 3 P6
rlabel metal1 -1713 880 -1706 881 5 P7
rlabel metal1 1360 -1665 1361 -1647 3 gnd
rlabel metal1 1545 -1697 1546 -1693 3 B3
rlabel metal1 1543 -1783 1544 -1779 3 B2
rlabel metal1 1546 -1869 1547 -1865 3 B1
rlabel metal1 1541 -2325 1542 -2321 3 B0
rlabel metal1 1583 -1651 1584 -1642 7 A0
rlabel metal1 1535 -1138 1535 -1134 3 B3
rlabel metal1 1537 -1224 1537 -1220 3 B2
rlabel metal1 1539 -1310 1539 -1306 3 B1
rlabel metal1 1538 -1396 1538 -1392 3 B0
rlabel metal1 425 -279 425 -275 3 B3
rlabel metal1 426 -365 426 -361 3 B2
rlabel metal1 427 -451 427 -447 3 B1
rlabel metal1 428 -537 428 -533 3 B0
rlabel metal1 -664 580 -664 584 3 B3
rlabel metal1 -663 494 -663 498 3 B2
rlabel metal1 -661 408 -661 412 3 B1
rlabel metal1 -662 322 -662 326 3 B0
rlabel metal1 -619 611 -619 615 3 A3
rlabel metal1 474 -245 474 -241 3 A2
rlabel metal1 1580 -1103 1580 -1099 3 A1
<< end >>
