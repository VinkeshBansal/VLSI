.INCLUDE 22nm_MGK.pm


*NAND GATE 

****Parameters**********
.PARAM Lmin=22n
.PARAM Wmin=22n
.PARAM XX=1
.PARAM tr=10p
.PARAM pvdd= 1

.temp 25

***Supply**************
vgndd gndd! 0 dc=0
vvddd vddd! 0 dc='pvdd'


****Capacitive load******


*MOSNAME drain gate source body type w l

****Net-list*************
.subckt adder nodeA nodeB nodeC nodesum nodecarry vddd! gndd!
Mn1	node11	nodeA	gndd!	gndd! 	nmos W={1*XX*Wmin} L={Lmin}
Mn2	node10	nodeA	gndd!	gndd! 	nmos W={1*XX*Wmin} L={Lmin}
Mn3	node10	nodeB	gndd!	gndd! 	nmos W={1*XX*Wmin} L={Lmin}
Mn4	node9	nodeC	gndd!	gndd! 	nmos W={1*XX*Wmin} L={Lmin}
Mn5	node9	nodeA	gndd!	gndd! 	nmos W={1*XX*Wmin} L={Lmin}
Mn6	node9	nodeB	gndd!	gndd! 	nmos W={1*XX*Wmin} L={Lmin}
Mn7	node8	nodeA	gndd!	gndd! 	nmos W={1*XX*Wmin} L={Lmin}
Mn8	node7	nodeB	node8	gndd! 	nmos W={1*XX*Wmin} L={Lmin}
Mn9	node6	nodeC	node7	gndd! 	nmos W={1*XX*Wmin} L={Lmin}
Mn10	node6	node12	node9	gndd! 	nmos W={1*XX*Wmin} L={Lmin}
Mn11	node12	nodeC	node10	gndd! 	nmos W={1*XX*Wmin} L={Lmin}
Mn12	node12	nodeB	node11	gndd! 	nmos W={1*XX*Wmin} L={Lmin}
Mp1	node1	nodeA	vddd!	vddd! 	pmos W={2*XX*Wmin} L={Lmin}
Mp2	node2	nodeA	vddd!	vddd! 	pmos W={2*XX*Wmin} L={Lmin}
Mp3	node2	nodeB	vddd!	vddd! 	pmos W={2*XX*Wmin} L={Lmin}
Mp4	node3	nodeC	vddd!	vddd! 	pmos W={2*XX*Wmin} L={Lmin}
Mp5	node3	nodeA	vddd!	vddd! 	pmos W={2*XX*Wmin} L={Lmin}
Mp6	node3	nodeB	vddd!	vddd! 	pmos W={2*XX*Wmin} L={Lmin}
Mp7	node4	nodeA	vddd!	vddd! 	pmos W={2*XX*Wmin} L={Lmin}
Mp8	node5	nodeB	node4	vddd! 	pmos W={2*XX*Wmin} L={Lmin}
Mp9	node6	nodeC	node5	vddd! 	pmos W={2*XX*Wmin} L={Lmin}
Mp10	node6	node12	node3	vddd! 	pmos W={2*XX*Wmin} L={Lmin}
Mp11	node12	nodeC	node2	vddd! 	pmos W={2*XX*Wmin} L={Lmin}
Mp12	node12	nodeB	node1	vddd! 	pmos W={2*XX*Wmin} L={Lmin}
Mp13    nodesum node6  vddd!   vddd!    pmos W={2*XX*Wmin} L={Lmin}
Mp14    nodecarry node12  vddd!   vddd!    pmos W={2*XX*Wmin} L={Lmin}
Mn13    nodesum node6  gndd!   gndd!    nmos W={1*XX*Wmin} L={Lmin}
Mn14    nodecarry node12  gndd!   gndd!    nmos W={1*XX*Wmin} L={Lmin}

.ends adder

.subckt and nodeA nodeB node6 vddd! gndd!
Mp1	node5	nodeA	vddd!	vddd! 	pmos W={2*XX*Wmin} L={Lmin}
Mp2	node5	nodeB	vddd! 	vddd! 	pmos W={2*XX*Wmin} L={Lmin} 
Mn1	node4	nodeA	gndd! 	gndd! 	nmos W={1*XX*Wmin} L={Lmin}
Mn2	node5	nodeB	node4 	gndd! 	nmos W={1*XX*Wmin} L={Lmin}
Mn3 node6   node5   gndd!   gndd!   nmos W={1*XX*Wmin} L={Lmin}
Mp3 node6   node5   vddd!   vddd!   pmos W={2*XX*Wmin} L={Lmin}  
.ends and


Xa1 nodeB3 nodeA3 nodeP vddd! gndd! and
Xa2 nodeB2 nodeA3 nodeO vddd! gndd! and
Xa3 nodeB3 nodeA2 nodeN vddd! gndd! and
Xa4 nodeB3 nodeA1 nodeM vddd! gndd! and
Xa5 nodeB1 nodeA3 nodeL vddd! gndd! and
Xa6 nodeB2 nodeA2 nodeK vddd! gndd! and
Xa7 nodeB1 nodeA2 nodeJ vddd! gndd! and
Xa8 nodeB0 nodeA3 nodeI vddd! gndd! and
Xa9 nodeB3 nodeA0 nodeH vddd! gndd! and 
Xa10 nodeB2 nodeA1 nodeG vddd! gndd! and
Xa11 nodeB1 nodeA1 nodeF vddd! gndd! and
Xa12 nodeB0 nodeA2 nodeE vddd! gndd! and
Xa13 nodeB2 nodeA0 nodeD vddd! gndd! and
Xa14 nodeB0 nodeA1 nodeC vddd! gndd! and
Xa15 nodeB1 nodeA0 nodeB vddd! gndd! and
Xa16 nodeB0 nodeA0 nodeP0 vddd! gndd! and

Xf1 nodeB nodeC 0 nodeP1 nodeha1c vddd! gndd! adder
Xf2 nodeE nodeF 0 nodeha2s nodeha2c vddd! gndd! adder
Xf3 nodeI nodeJ 0 nodeha3s nodeha3c vddd! gndd! adder
Xf4 nodeN nodeO nodefa7c nodefa4s nodefa4c vddd! gndd! adder
Xf5 nodeD nodeha1c nodeha2s nodeP2 nodefa5c vddd! gndd! adder
Xf6 nodeG nodeha2c nodeha3s nodefa6s nodefa6c vddd! gndd! adder
Xf7 nodeK nodeL nodeha3c nodefa7s nodefa7c vddd! gndd! adder
Xf8 nodeP nodefa4c nodefa12c nodeP6 nodeC5 vddd! gndd! adder
Xf9 nodefa5c nodefa6s nodeH nodeP3 nodefa9c vddd! gndd! adder
Xf10 nodefa9c nodefa11s 0 nodeP4 nodeha10c vddd! gndd! adder
Xf11 nodefa7s nodefa6c nodeM nodefa11s nodefa11c vddd! gndd! adder
Xf12 nodeha10c nodefa11c nodefa4s nodeP5 nodefa12c vddd! gndd! adder


Cout  nodeP0 0 2f
Cout  nodeP1 0 2f
Cout  nodeP2 0 2f
Cout  nodeP3 0 2f
Cout  nodeP4 0 2f
Cout  nodeP5 0 2f
Cout  nodeP6 0 2f
Cout  nodeC5 0 2f


*******input**********




VinA0 nodeA0 0 pulse 0 1 0 100p 100p 50n 100n
VinA1 nodeA1 0 pulse 0 1 0 100p 100p 100n 200n
VinA2 nodeA2 0 pulse 0 1 0 100p 100p 200n 400n
VinA3 nodeA3 0 pulse 0 1 0 100p 100p 400n 800n
VinB0 nodeB0 0 pulse 0 1 0 100p 100p 800n 1600n
VinB1 nodeB1 0 pulse 0 1 0 100p 100p 1600n 3200n
VinB2 nodeB2 0 pulse 0 1 0 100p 100p 3200n 6400n
VinB3 nodeB3 0 pulse 0 1 0 100p 100p 6400n 12800n
* analysis mode
.TRAN 1n 12800n




*measure
* .meas tran delay_LHB trig V(nodeB) val=0.5 fall=2 targ V(node5) val=0.5 rise=3
* .meas tran delay_HLA trig V(nodeA) val=0.5 rise=2 targ V(node5) val=0.5 fall=2
* .meas tran delay_LHA trig V(nodeA) val=0.5 fall=2 targ V(node5) val=0.5 rise=2
* .meas tran delay_HLB trig V(nodeB) val=0.5 rise=1 targ V(node5) val=0.5 fall=1

 
.control
run
plot nodeP0+14 nodeP1+12 nodeP2+10 nodeP3+8 nodeP4+6 nodeP5+4 nodeP6+2 nodeC5 nodeA3-2 nodeA2-4 nodeA1-6 nodeA0-8 nodeB3-10 nodeB2-12 nodeB1-14 nodeB0-16
.endc

.end
